`timescale  1ns/1ns

module tb_fifo_8to3();
reg		clock,rst_n,r_en,w_en;
reg	[7:0]	in_data;
wire	[2:0]	out_data;
wire		full,empty,half_full,overflow;

reg     [2:0]   out_golden_data;
reg		out_golden_full, out_golden_empty, out_golden_half_full, out_golden_overflow;

integer i;

//used reg to simulate queue
reg [127:0] data_stored;
reg [7:0] space_avail;
reg [6:0] head_fifo_ptr;
reg [6:0] tail_fifo_ptr;

//GENERAL RULES FOR TESTBENCH:

//ON THE NEGEDGE OF CLOCK SIGNAL, THE INPUT SIGNAL FOR THE DUT MODULE AND THE OUTPUT GOLDEN SIGNALS GENERATED BY THE OUTPUT GOLDEN MODEL ARE GENERATED AT THE SAME TIME
//==============================
//ONE PERIOD AHEAD OF THE POSEDGE, WHEN THE DUT PRODUCED THE OUTPUT SIGNALS
//===============================
//ON THE FOLLOWING NEGEDGE, COMPARE THE DUT OUTPUT WITH THE GOLDEN OUTPUT
//========================
//A TEST IS DONE ONCE FOR THIS INPUT

//READ AND WRITE AT THE SAME TIME IS NOT TESTED

//queue pop function
//this chunk of code is meant to be serially conducted
//so written in C style
task read;
	input r_en;
	output [2:0] out_golden_data;
	output out_golden_full;
	output out_golden_empty;
	output out_golden_half_full;
	output out_golden_overflow;

	if(r_en) begin
		if(space_avail == 8'd128) begin
			$display("CAN'T READ WHEN FIFO IS EMPTY\n");
			$stop;
		end
		else if(space_avail == 8'd127) begin
			$display("CAN'T READ WHEN FIFO IS EMPTY\n");
			$stop;
		end
		else if(space_avail == 8'd126) begin
			$display("CAN'T READ WHEN FIFO IS EMPTY\n");
			$stop;
		end
		else begin
			if(head_fifo_ptr == 7'd126) begin
				space_avail = space_avail + 3;
				out_golden_data = {data_stored[0] ,data_stored[127:126]};
				head_fifo_ptr = 6'd1;
			end

			else if(head_fifo_ptr == 7'd127) begin
				space_avail = space_avail + 3;
				out_golden_data = {data_stored[1:0], data_stored[127]};
				head_fifo_ptr = 6'd2;
			end

			else begin
				space_avail = space_avail + 3;
				out_golden_data = {data_stored[head_fifo_ptr[6:0] +: 3]};
				//The problem is that in Verilog you can't have two variable expressions in a range, even if they evaluate to a constant difference.
				//An error occur if change to [head_fifo_ptr[5:0] + 3 : head_fifo_ptr[5:0]].
				head_fifo_ptr = head_fifo_ptr + 3;
			end

			if(space_avail == 7'd64) 
				out_golden_half_full = 1'b1;
			else
				out_golden_half_full = 1'b0;

			if(space_avail >= 7'd126)
				out_golden_empty = 1'b1;
			else
				out_golden_empty = 1'b0;

			out_golden_full = 1'b0;
			out_golden_overflow = 1'b0;
		end
	end


endtask

//queue push function
task write;
	input w_en;
	input [7:0] in_data;
	output out_golden_full;
	output out_golden_empty;
	output out_golden_half_full;
	output out_golden_overflow;

	if(w_en) begin
		if(space_avail < 7'd8) begin
			out_golden_overflow = 1'b1;
			out_golden_full = 1'b1;
			out_golden_empty = 1'b0;
			out_golden_half_full = 1'b0;
			$display("CAN'T WRITE WHEN FIFO IS FULL, OVERFLOW\n");
		end
		else begin
			data_stored[tail_fifo_ptr[6:0] +: 8] = in_data;
			tail_fifo_ptr = tail_fifo_ptr + 8;
			space_avail = space_avail - 8;
		
		
			if(space_avail == 7'd64) 
				out_golden_half_full = 1'b1;
			else
				out_golden_half_full = 1'b0;

			if(space_avail < 7'd8)
				out_golden_full = 1'b1;
			else
				out_golden_full = 1'b0;
			out_golden_empty = 1'b0;
			out_golden_overflow = 1'b0;
		end
	end

	else
		out_golden_overflow = 1'b0;

endtask


fifo	FIFO(    
		.clk(clock),
		 .rst_n(rst_n),
		 .w_en(w_en),
		 .data_w(in_data),
		 .r_en(r_en),
		 .data_r(out_data),
		 .empty(empty),
		 .full(full),
		 .half_full(half_full),
		 .overflow(overflow));

initial
begin
    in_data=0;
	r_en=0;
	w_en=0;
	clock=1;
	rst_n=0;
	i=1;

	space_avail = 8'd128;
	head_fifo_ptr = 7'd0;
	tail_fifo_ptr = 7'd0;

	//initialize the out_golden_signals
	out_golden_empty = 1'b1;
	out_golden_full = 1'b0;
	out_golden_half_full = 1'b0;
	out_golden_overflow = 1'b0;

	#25 rst_n=1;
	$display("\n\ninitial done\n\n");
	if({empty,half_full,full,overflow}!={out_golden_empty, out_golden_half_full, out_golden_full, out_golden_overflow})
	begin
		$display("\nerror at time %0t:",$time);
		$display("after reset,status not asserted\n");
		$display("empty = %b full = %b half_full = %b overflow = %b\n",empty,full,half_full,overflow);
		$stop;
	end
	else
	begin
		$display("initial status right\nempty = %b full = %b half_full = %b overflow = %b\n",empty,full,half_full,overflow);
	end
   #25;


	//causing half_full
	for (i=1;i<9;i=i+1)
	begin
	   @(negedge clock) w_en=1; in_data=i; write(w_en, in_data, out_golden_full, out_golden_empty, out_golden_half_full, out_golden_overflow);
		$display("storing %d  w_en=%d r_en=%d\n",i,w_en,r_en);
	end
	@(negedge clock) w_en=0;
	#10;
	if({empty,half_full,full,overflow}!={out_golden_empty, out_golden_half_full, out_golden_full, out_golden_overflow})
	begin
		$display("\nerror at time %0t:",$time);
		$display("half_full\n");
		$display("empty = %b full = %b half_full = %b overflow = %b\n",empty,full,half_full,overflow);
		$stop;
	end
	else
	begin
		$display("half_full status right\nempty = %b full = %b half_full = %b overflow = %b\n",empty,full,half_full,overflow);
	end


	//causing full
	for (i=9;i<17;i=i+1)
	begin
	   @(negedge clock) w_en=1; in_data=i; write(w_en, in_data, out_golden_full, out_golden_empty, out_golden_half_full, out_golden_overflow);
		$display("storing %d  w_en=%d r_en=%d\n",i,w_en,r_en);
	end
	@(negedge clock) w_en=0;
	#25;
	if({empty,half_full,full,overflow}!={out_golden_empty, out_golden_half_full, out_golden_full, out_golden_overflow})
	begin
		$display("\nerror at time %0t:",$time);
		$display("full\n");
		$display("empty = %b full = %b half_full = %b overflow = %b\n",empty,full,half_full,overflow);
		$stop;
	end
	else
	begin
		$display("full status right\nempty = %b full = %b half_full = %b overflow = %b\n",empty,full,half_full,overflow);
	end

	//causing overflow
	begin
	   @(negedge clock) w_en=1;in_data = 99; write(w_en, in_data, out_golden_full, out_golden_empty, out_golden_half_full, out_golden_overflow);
		$display("storing %d  w_en=%d r_en=%d\n",i,w_en,r_en);
	end
	#25;
	if({empty,half_full,full,overflow}!={out_golden_empty, out_golden_half_full, out_golden_full, out_golden_overflow})
	begin
		$display("\nerror at time %0t:",$time);
		$display("overflow\n");
		$display("empty = %b full = %b half_full = %b overflow = %b\n",empty,full,half_full,overflow);
		$stop;
	end
	else
	begin
		$display("overflow status right\nempty = %b full = %b half_full = %b overflow = %b\n",empty,full,half_full,overflow);
	end
	//these nums r in fifo 1~16
	//starting to read nums
	//@(negedge clock) w_en=0;r_en=1; denote this line because the input and the golden model need change at the same time
	for (i=1;i<5;i=i+1)
	begin
	   @(negedge clock) r_en = (i == 4) ? 0 : 1; w_en = 0;
	   	read(r_en, out_golden_data, out_golden_full, out_golden_empty, out_golden_half_full, out_golden_overflow);
		#7;
		//can't be #5, dut module has delay time after the posedge of clk to produce the output  
		$display("Iteration %d, r_en = %d, reading data %d, your data %d\n",i,r_en,out_golden_data,out_data);
		//wait for the output of dut model and then compare
		if(out_data!=out_golden_data)
		begin
			$display("expected data %d\n your data %d",out_golden_data,out_data);
		$stop;
		end
	end

	#25;
	if({empty,half_full,full,overflow}!={out_golden_empty, out_golden_half_full, out_golden_full, out_golden_overflow})
	begin
		$display("\nerror at time %0t:",$time);
		$display("empty = %b full = %b half_full = %b overflow = %b\n",empty,full,half_full,overflow);
		$stop;
	end
	else
	begin
		$display("after reading 4 data, right, empty = %b full = %b half_full = %b overflow = %b\n",empty,full,half_full,overflow);
	end
	
	@(negedge clock) r_en=0;
	#25;
	for (i=1;i<5;i=i+1)  
	begin
	   @(negedge clock) w_en=1;in_data=i; write(w_en, in_data, out_golden_full, out_golden_empty, out_golden_half_full, out_golden_overflow);
		$display("storing %d again  w_en=%d r_en=%d\n",i,w_en,r_en);
	end

	#25;
	if({empty,half_full,full,overflow}!={out_golden_empty, out_golden_half_full, out_golden_full, out_golden_overflow})
	begin
		$display("\nerror at time %0t:",$time);
		$display("overflow\n");
		$display("empty = %b full = %b half_full = %b overflow = %b\n",empty,full,half_full,overflow);
		$stop;
	end
	else
	begin
		$display("overflow status right\nempty = %b full = %b half_full = %b overflow = %b\n",empty,full,half_full,overflow);
	end

	//read fifo all out, there are 41 3-bit data in the fifo
	//@(negedge clock) w_en=0; r_en=1;	
	//i < 43 get "done without error"
	//i < 44 get "CAN'T READ WHEN FIFO IS EMPTY"
	for (i=1;i<44;i=i+1)
	begin
	   @(negedge clock) r_en = (i == 44) ? 0 : 1; w_en = 0;
		read(r_en, out_golden_data, out_golden_full, out_golden_empty, out_golden_half_full, out_golden_overflow);
		#7;
		$display("reading data %d  actually get %d\n",out_golden_data,out_data);		
		if(out_data!=out_golden_data)
		begin
			$display("date stored in %d maybe wrong\n",out_data);
			$stop;
		end	
	end

	#25;
	if({empty,half_full,full,overflow}!={out_golden_empty, out_golden_half_full, out_golden_full, out_golden_overflow})
	begin
		$display("\nerror at time %0t:",$time);
		$display("empty = %b full = %b half_full = %b overflow = %b\n",empty,full,half_full,overflow);
		$stop;
	end
	else
	begin
		$display("********************\ndone, without error\n********************\n");
		$stop;
	end
	


end

always #5 clock = ~clock;

endmodule